module div (
    input [7:0] n1,
    input [7:0] n2,
    output [7:0] div
);
    assign  div=n1/n2;

endmodule