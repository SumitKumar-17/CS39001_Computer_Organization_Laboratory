module mult (
    input [7:0] n1,
    input [7:0] n2,
    output [7:0] mult
);
    assign  mult=n1*n2;

endmodule