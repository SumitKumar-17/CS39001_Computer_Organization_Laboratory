`timescale 1ns / 1ps

module outeqinp(
     input [31:0] a,
     output [31:0] out
);
    assign out=a;
endmodule
